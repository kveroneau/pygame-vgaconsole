� �  �QBASIC   EXE            194,309 21-12-2014 22:54                                QBASIC   HLP            130,881 21-12-2014 22:54                                    2 File(s)           325,190 Bytes.                                              2 Dir(s)        262,111,744 Bytes free.                                                                                                                     C:\QBASIC>QBASIC.EXE                                                                                                                                            Type EXIT to return to QBasic                                                   ����������������������������������������������������������������������          � Welcome to DOSBox v0.74                                            �          �                                                                    �          � For a short introduction for new users type: INTRO                 �          � For supported shell commands type: HELP                            �          �                                                                    �          � To adjust the emulated CPU speed, use ctrl-F11 and ctrl-F12.       �          � To activate the keymapper ctrl-F1.                                 �          � For more information read the README file in the DOSBox directory. �          �                                                                    �          � HAVE FUN!                                                          �          � The DOSBox Team http://www.dosbox.com                              �          ����������������������������������������������������������������������          C:\QBASIC>exit                                                                                                                                                                                                                                                                                                                  